-------------------------------------------------------------------------------
--
-- Title       : ALU Register Decoder
-- Author      : Matthew Champagne
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- Generated   : Wed Nov 26 18:25:15 2021
--
-------------------------------------------------------------------------------
--
-- Description : Takes all the inputs generated by the instruction and chooses
-- which fields go into the ALU.
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;


entity ALURegisterDecoder is 
	port(
		--Input
		cop : in std_logic_vector(4 downto 0);
		valueA : in std_logic_vector(127 downto 0);
		valueB : in std_logic_vector(127 downto 0);
		valueC : in std_logic_vector(127 downto 0);
		loadIndex : in std_logic_vector(2 downto 0);
		immediate : in std_logic_vector(15 downto 0);
		forward : in std_logic_vector(2 downto 0);
		forwardValue : in std_logic_vector(127 downto 0); 
		
		--Output
		rs1 : out std_logic_vector(127 downto 0);
		rs2 : out std_logic_vector(127 downto 0);
		rs3 : out std_logic_vector(127 downto 0)
	);
end ALURegisterDecoder;		


architecture behavioral of ALURegisterDecoder is
	begin										 							  
	
		decode : process(cop, valueA, valueB, valueC, loadIndex, immediate, forward, forwardValue)
			begin					   		
				rs1 <= valueA;
				rs2 <= valueB;
				rs3 <= valueC;
					
				if(forward(0 downto 0) = "1") then
					rs1 <= forwardValue;
					
				end if;
					
				if(forward(1 downto 1) = "1") then
					rs2 <= forwardValue;
					
				end if;
				
				if(forward(2 downto 2) = "1") then
					rs3 <= forwardValue;
					
				end if;
					
					
				--Special case loadImmediate
				if(to_integer(unsigned(cop(4 downto 0))) = 0) then
					rs1 <= std_logic_vector(to_unsigned(0, 128)); --clears output to all zeros
					rs1(15 downto 0) <= immediate;

					rs2 <= std_logic_vector(to_unsigned(0, 128)); --clears output to all zeros
					rs2(2 downto 0) <= loadIndex;
					
				--Special case Shift Left Halfword Immediate
				elsif(to_integer(unsigned(cop(4 downto 0))) = 21) then
					rs1 <= valueA;	
					
					rs2 <= std_logic_vector(to_unsigned(0, 128)); --clears output to all zeros
					rs2(4 downto 0) <= immediate(9 downto 5);
					
				end if;
		end process;
end behavioral;